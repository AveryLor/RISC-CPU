module control_unit(SW, LEDR, KEY, HEX0, HEX1);
  // Hardware I/O
  input [9:0] SW;
  input [2:0] KEY;
  output [9:0] LEDR;
  output [6:0] HEX0;
  output [6:0] HEX1;

  // Necessary values
  wire [7:0] instruction_state = SW[7:0];

  // Clock pulse and reset
  wire clock_pulse = ~KEY[0];
  wire resetn = KEY[1];
  wire stall = ~KEY[2]; // This will be changed later. It is kept just for testing the module.

  // Registers
  wire [31:0] IR; // Special purpose
  /* Should add 16-bit pc register when program counter is implemented. */
  
  // Pipeline registers
  wire [7:0] if_id_reg;
 
  wire id_ex_regwrite;
  wire id_ex_reg_mode;
  wire [2:0] id_ex_reg_opcode;
  wire [31:0] id_ex_reg_val1;
  wire [31:0] id_ex_reg_val2;
  wire [1:0] id_ex_reg_wb_enc; 
  
  wire ex_mem_regwrite;
  wire [31:0] ex_mem_reg_arithmetic_result;
  wire [1:0] ex_mem_reg_wb_enc;

  wire mem_wb_regwrite;
  wire [1:0] mem_wb_reg_wb_enc;
  wire [31:0] mem_wb_reg_arithmetic_result;

  // Register file conntrol
  wire we;
  wire [31:0] wdata; 
  wire [1:0] r_write_enc;

  wire [1:0] r_enc_0;
  wire [1:0] r_enc_1;

  wire [31:0] rf_out_val1;
  wire [31:0] rf_out_val2;

  wire [31:0] R0_val;
  wire [31:0] R1_val;

  reg_file reg_file_inst(
      .clk(clock_pulse),
      .resetn(resetn),

      .we(we),

      .r_enc_0(r_enc_0),
      .r_enc_1(r_enc_1),

      .r_write_enc(r_write_enc),

      .reg_out_0(rf_out_val1),
      .reg_out_1(rf_out_val2),

      .wdata(wdata),

      .R0_val(R0_val),
      .R1_val(R1_val)
  );

  // Hex display for register file
  display_hex display_hex_inst0(R0_val, HEX0);
  display_hex display_hex_inst1(R1_val, HEX1);

  // ALU Control 
  wire [2:0] alu_opcode;
  wire [31:0] alu_reg_val1;
  wire [31:0] alu_reg_val2;
  wire [31:0] alu_result; 

  // ALU instantiation
  ALU alu_inst(
    .opcode(alu_opcode),
    .arithmetic_result(alu_result), 
    .register_value_1(alu_reg_val1),
    .register_value_2(alu_reg_val2)
  );
  
  instr_fetch instr_fetch_inst(
      .clk(clock_pulse),
      .stall(stall)
	  .pc(), // add 16-bit program counter here
      .switches_state(instruction_state),
      .if_id_reg(if_id_reg)
  );

  instr_decode instr_decode_inst(
      .clk(clock_pulse),
      .stall(stall),

      .rf_enc_0(r_enc_0),
      .rf_enc_1(r_enc_1),

      .rf_out_val1(rf_out_val1),
      .rf_out_val2(rf_out_val2),

      .if_id_reg(if_id_reg), 

      .id_ex_reg_val1(id_ex_reg_val1),
      .id_ex_reg_val2(id_ex_reg_val2), 
      .id_ex_reg_mode(id_ex_reg_mode),
      .id_ex_reg_opcode(id_ex_reg_opcode),
      .id_ex_reg_wb_enc(id_ex_reg_wb_enc),
      .id_ex_regwrite(id_ex_regwrite)
  );

  instr_execute instr_execute_inst(
      .clk(clock_pulse),

      .alu_opcode(alu_opcode),
      .alu_reg_val1(alu_reg_val1),
      .alu_reg_val2(alu_reg_val2),
      .alu_result(alu_result),
      
      .id_ex_reg_opcode(id_ex_reg_opcode),
      .id_ex_reg_val1(id_ex_reg_val1),
      .id_ex_reg_val2(id_ex_reg_val2),
      .id_ex_regwrite(id_ex_regwrite),
      .id_ex_reg_wb_enc(id_ex_reg_wb_enc),

      .ex_mem_reg_wb_enc(ex_mem_reg_wb_enc),
      .ex_mem_regwrite(ex_mem_regwrite),
      .ex_mem_reg_arithmetic_result(ex_mem_reg_arithmetic_result)
  ); 
  
  instr_mem instr_mem_inst(
      .clk(clock_pulse),

      .ex_mem_regwrite(ex_mem_regwrite),
      .ex_mem_reg_wb_enc(ex_mem_reg_wb_enc),
      .ex_mem_reg_arithmetic_result(ex_mem_reg_arithmetic_result),

      .mem_wb_reg_wb_enc(mem_wb_reg_wb_enc),
      .mem_wb_reg_arithmetic_result(mem_wb_reg_arithmetic_result),
      .mem_wb_regwrite(mem_wb_regwrite)

  );

  instr_wb instr_wb_inst(
      .clk(clock_pulse),

      .mem_wb_regwrite(mem_wb_regwrite),
      .mem_wb_reg_wb_enc(mem_wb_reg_wb_enc),
      .mem_wb_reg_arithmetic_result(mem_wb_reg_arithmetic_result),

      .rf_we(we),
      .rf_w_enc(r_write_enc),
      .rf_wdata(wdata)
  );
  
  // Testing decode: 
  assign LEDR[2:0] = ex_mem_reg_arithmetic_result;
  assign LEDR[8:7] = mem_wb_reg_wb_enc;
  assign LEDR[9] = mem_wb_regwrite;
  //assign LEDR[9:7] = if_id_reg[6:4];
  //assign LEDR[6:4] = id_ex_reg_opcode; 
  //assign LEDR[3:2] = ex_mem_regwrite;
  //assign LEDR[1:0] = mem_wb_regwrite;
endmodule

// Register file module 
module reg_file(clk, resetn, we, r_enc_0, r_enc_1, r_write_enc, reg_out_0, reg_out_1, wdata, R0_val, R1_val, register_output); 
  input we; // Indicates if we are doing a write (write enable)
  input clk;
  input resetn;

  input [1:0] r_enc_0; // Register encodings 
  input [1:0] r_enc_1; 
  input [1:0] r_write_enc;
  input [31:0] wdata;

  output [31:0] R0_val;
  output [31:0] R1_val;
  
  output [31:0] register_output[7:0];

  output reg [31:0] reg_out_0;
  output reg [31:0] reg_out_1;
  
  // The actual registers =)
  reg [31:0] R0;
  reg [31:0] R1;

  // Reading registers
  // We use blocking assignments here because it behaves a little better in simulation.
  always @ (*) begin
    reg_out_0 = (r_enc_0 == 2'b00) ? R0 : R1;
    reg_out_1 = (r_enc_1 == 2'b00) ? R0 : R1;
  end
  
  // Writing to registers.
  always @ (posedge clk or negedge resetn) begin
    if (!resetn) begin
      R0 <= 32'd3;
      R1 <= 32'd3;
    end
    else if (we) begin
      if (r_write_enc == 2'b00) R0 <= wdata;
      else R1 <= wdata; 
    end
  end

  assign register_output[0] = R0;
  assign register_output[1] = R1;
  assign register_output[2] = R2; 
  assign register_output[3] = R3;
  assign register_output[4] = R4;
  assign register_output[5] = R5;
  assign register_output[6] = R6;
  assign register_output[7] = R7;

endmodule


// ALU Module
module ALU(opcode, arithmetic_result, register_value_1, register_value_2);
  parameter [2:0] ADD = 3'b001,
                  INC = 3'b011;

  input [2:0] opcode;
  input [31:0] register_value_1;
  input [31:0] register_value_2;
  
  output reg [31:0] arithmetic_result;
  always @ (*) begin
    case (opcode) 
      ADD: arithmetic_result = register_value_1 + register_value_2; 
      INC: arithmetic_result = register_value_1 + 1; 
      default: arithmetic_result = 32'b0;
    endcase
  end
endmodule


module instr_fetch(clk, stall, pc, switches_state, if_id_reg);
  input clk;
  input stall;
  input [15:0] pc;				// program counter (new)
  input [7:0] switches_state; 	// no longer used
  output [31:0] if_id_reg;		// changed to 32 bits. instead of a reg, this is now a wire to a BRAM DataOut reg.
  
  /* START OF NEW ADDITIONS */
  // This module will be defined by quartus. 
  // In Quartus, name the BRAM instr_rom, set width = 32, depth = 65536, use a single clock, and initialize it with a .mif.
  
  instr_rom instr_rom(
	.address(pc),
	.clock(clk),
	.data()
	.wren(0),
	.q(if_id_reg);

	input	[15:0]  address;
	input	clock;
	input	[7:0]  data;
	input	wren;
	output	[7:0]  q;
  );
  
  /* END OF NEW ADDITIONS */

  // If you want to stall here, just keep the program counter static instead.
  /*
  always @ (posedge clk) begin 
    if (stall == 0) if_id_reg <= switches_state;
    else if_id_reg <= if_id_reg;
  end
  */
endmodule

module instr_decode(clk, stall, rf_enc_0, rf_enc_1, rf_out_val1, rf_out_val2, if_id_reg, id_ex_reg_val1, id_ex_reg_val2, id_ex_reg_mode, id_ex_reg_opcode, id_ex_reg_wb_enc, id_ex_regwrite);
  input clk;
  input stall;
  input [7:0] if_id_reg;

  
  output reg id_ex_reg_mode;
  output reg [2:0] id_ex_reg_opcode;
  output reg [1:0] id_ex_reg_wb_enc;
  output reg id_ex_regwrite;

  output reg [31:0] id_ex_reg_val1;
  output reg [31:0] id_ex_reg_val2;

  // Register file control
  output [1:0] rf_enc_0;
  output [1:0] rf_enc_1;

  input [31:0] rf_out_val1;
  input [31:0] rf_out_val2;
  
  // Must be purely combinational to get timing right.
  assign rf_enc_0 = if_id_reg[3:2];
  assign rf_enc_1 = if_id_reg[1:0];
  
  // values will be given by the register file once it is instantiated.
  always @ (posedge clk) begin
    if (!stall) begin
      id_ex_reg_mode <= if_id_reg[7];
      id_ex_reg_opcode <= if_id_reg[6:4];
      id_ex_reg_wb_enc <= if_id_reg[3:2];

      id_ex_reg_val1 <= rf_out_val1;
      id_ex_reg_val2 <= rf_out_val2;

      if (if_id_reg[6:4] != 3'b000) id_ex_regwrite <= 1;
      else id_ex_regwrite <= 0;
    end
  end
endmodule

module instr_execute(clk, alu_opcode, alu_reg_val1, alu_reg_val2, alu_result, id_ex_reg_opcode, id_ex_reg_val1, id_ex_reg_val2, id_ex_regwrite, id_ex_reg_wb_enc, ex_mem_reg_wb_enc, ex_mem_regwrite, ex_mem_reg_arithmetic_result);
  input clk;
  
  // From ID/EX pipeline
  input        id_ex_regwrite;
  input [1:0]  id_ex_reg_wb_enc;
  input [2:0]  id_ex_reg_opcode;
  input [31:0] id_ex_reg_val1;
  input [31:0] id_ex_reg_val2;

  // EX/MEM pipeline registers
  output reg [1:0] ex_mem_reg_wb_enc;
  output reg ex_mem_regwrite;
  output reg [31:0] ex_mem_reg_arithmetic_result;
  
  // To ALU (combinational - wires)  
  output [2:0] alu_opcode;

  output [31:0] alu_reg_val1;
  output [31:0] alu_reg_val2;
  
  // ALU output
  input [31:0] alu_result;
  
  assign alu_opcode = id_ex_reg_opcode;
  assign alu_reg_val1 = id_ex_reg_val1;
  assign alu_reg_val2 = id_ex_reg_val2;

  always @ (posedge clk) begin
    ex_mem_reg_wb_enc <= id_ex_reg_wb_enc;
    ex_mem_regwrite <= id_ex_regwrite;
    ex_mem_reg_arithmetic_result <= alu_result;
  end
endmodule

module instr_mem(clk, ex_mem_regwrite, ex_mem_reg_wb_enc, ex_mem_reg_arithmetic_result, mem_wb_reg_wb_enc, mem_wb_reg_arithmetic_result, mem_wb_regwrite);
  input clk;
  input [1:0] ex_mem_reg_wb_enc;
  input [31:0] ex_mem_reg_arithmetic_result;
  input ex_mem_regwrite;
  
  output reg [1:0] mem_wb_reg_wb_enc;
  output reg [31:0] mem_wb_reg_arithmetic_result;
  output reg mem_wb_regwrite;
  
  always @ (posedge clk) begin
    mem_wb_reg_wb_enc <= ex_mem_reg_wb_enc;
    mem_wb_reg_arithmetic_result <= ex_mem_reg_arithmetic_result;
    mem_wb_regwrite <= ex_mem_regwrite;
  end
endmodule


module instr_wb(clk, mem_wb_regwrite, mem_wb_reg_wb_enc, mem_wb_reg_arithmetic_result, rf_we, rf_w_enc, rf_wdata); 
  input clk;

  input mem_wb_regwrite;
  input [1:0] mem_wb_reg_wb_enc;
  input [31:0] mem_wb_reg_arithmetic_result;

  output reg rf_we;
  output reg [1:0] rf_w_enc; 
  output reg [31:0] rf_wdata;

  always @ (posedge clk) begin
    rf_we <= mem_wb_regwrite;
    rf_w_enc <= mem_wb_reg_wb_enc; 
    rf_wdata <= mem_wb_reg_arithmetic_result;
  end
endmodule

/* Hex display module for displaying first few bytes of the registers on the hex displays*/
module display_hex(input [3:0] dig, output [6:0] HEX);
    reg [6:0] temp;
    assign HEX = temp;   // connect internal signal to output

    always @ (*) begin
        if (dig == 4'h0)
            temp = 7'b1000000;  // 0
        else if (dig == 4'h1)
            temp = 7'b1111001;  // 1
        else if (dig == 4'h2)
            temp = 7'b0100100;  // 2
        else if (dig == 4'h3)
            temp = 7'b0110000;  // 3
        else if (dig == 4'h4)
            temp = 7'b0011001;  // 4
        else if (dig == 4'h5)
            temp = 7'b0010010;  // 5
        else if (dig == 4'h6)
            temp = 7'b0000010;  // 6
        else if (dig == 4'h7)
            temp = 7'b1111000;  // 7
        else if (dig == 4'h8)
            temp = 7'b0000000;  // 8
        else if (dig == 4'h9)
            temp = 7'b0010000;  // 9
        else if (dig == 4'hA)
            temp = 7'b0001000;  // A
        else if (dig == 4'hB)
            temp = 7'b0000011;  // b
        else if (dig == 4'hC)
            temp = 7'b1000110;  // C
        else if (dig == 4'hD)
            temp = 7'b0100001;  // d
        else if (dig == 4'hE)
            temp = 7'b0000110;  // E
        else if (dig == 4'hF)
            temp = 7'b0001110;  // F
        else
            temp = 7'b1111111;  // display off (invalid input)
    end
endmodule
